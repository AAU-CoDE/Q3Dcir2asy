* BEGIN ANSOFT HEADER
* node 1    Net1:L1B
* node 2    Net2:L2B
* node 3    Net1:L1A
* node 4    Net2:L2A
*  Project: Q3Dcir2asy
*   Design: Q3DDesign1
*   Format: Ansys Nexxim
*   Topckt: parallel_conductors
*  Creator: Ansys Electronics Desktop 2024.2.0
*     Date: Wed Oct 02 13:20:13 2024
* END ANSOFT HEADER

.subckt parallel_conductors 1 2 3 4
XZhalf1 1 2 5 6 parallel_conductors_half
XY1 5 6 parallel_conductors_parlel
XZhalf2 5 6 3 4 parallel_conductors_half

.subckt parallel_conductors_half 1 2 3 4
L1 1 3 2.56779523113e-10
L2 2 4 2.568020091e-10
K1_2 L1 L2 0.295133
.ends parallel_conductors_half

.subckt parallel_conductors_parlel 1 2
.ends parallel_conductors_parlel

.ends parallel_conductors
